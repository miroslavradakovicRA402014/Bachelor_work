----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    14:47:40 04/13/2018 
-- Design Name: 
-- Module Name:    uart - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity uart is
    Port ( iCLK        		 : in   STD_LOGIC;
           inRST       		 : in   STD_LOGIC;
           iRX         		 : in   STD_LOGIC;
           iUART_RD    		 : in   STD_LOGIC;
           oUART_EMPTY      : out  STD_LOGIC;
           oUART_DATA       : out  STD_LOGIC_VECTOR (7 downto 0));
end uart;

architecture Behavioral of uart is

begin


end Behavioral;

